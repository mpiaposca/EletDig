library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package myDef is
  constant n:integer:=4;
end package myDef;
